module cornigera (
  input logic clk,
  address 
  datain
  dataout
);
 decode unit
 alu
 register_file
 load_unit
 store_unit
endmodule
