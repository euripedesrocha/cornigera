import cornigera_pkg::*;

module registers (
  input logic clk,
  input RegisterName write_to,
  input RegisterName read_from,
  input logic write_data,
  output logic read_date
);
endmodule
