package cornigera_pkg;
  typedef enum logic [4:0]{R0} RegisterName; 
endpackage
